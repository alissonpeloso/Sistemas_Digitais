module bc(
    
)